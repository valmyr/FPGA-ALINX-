module segment7(input [3:0] in, output [6:0] d);
	assign d  = (in == 0) ? 7'b0000001 :
		         (in == 1) ? 7'b1001111 :
					(in == 2) ? 7'b0010010 :
					(in == 3) ? 7'b0000110 :
					(in == 4) ? 7'b1001100 :
					(in == 5) ? 7'b0100100 :
					(in == 6) ? 7'b0100000 :
					(in == 7) ? 7'b0001111 :
					(in == 8) ? 7'b0000000 : 
					(in == 9) ? 7'b0000100 : 7'b1111111;
endmodule
